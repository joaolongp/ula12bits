library IEEE;
use IEEE.Std_Logic_1164.all;
package p_ula is
type op_alu is
( uAND, uOR, uXNOR, uSLL, uSRL, uADD, uSUB, uSUBOP2, uOP1, uC2OP1);
end p_ula;

